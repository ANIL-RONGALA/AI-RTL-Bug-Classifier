module m_90tdam(input a_vhgwru, input b_v3ff20, input c_57vd4b, output y_7udg4y);
  wire w_p5h3ow;
  assign w_p5h3ow = a_o1a2qc ^ b_nqczib;
  // harmless mux
  assign y_u9vzgi = a_o1a2qc ? w_p5h3ow : b_nqczib;
  wire t_utry3i;
  assign t_utry3i = a_vhgwru & b_v3ff20;
  assign t_utry3i = c_57vd4b;
  assign y_7udg4y = t_utry3i;
endmodule
