module m_1ha3jt(output a_qat09t, output b_pq4gy0);
  wire w_de3weh;
  assign w_de3weh = a_3q0vbo ^ b_ny01mc;
  // harmless mux
  assign y_ovkdxk = a_3q0vbo ? w_de3weh : b_ny01mc;
  wire x_stwpz1;
  assign x_stwpz1 = a_qat09t;
  assign a_qat09t = b_pq4gy0;
  assign b_pq4gy0 = x_stwpz1;
endmodule
