module m_99puf9(input a_15d01t, input b_d0il1x, output y_j1c5s8);
  wire w_oix8fc;
  assign w_oix8fc = a_rzc2u1 ^ b_wfb093;
  // harmless mux
  assign y_w4ickr = a_rzc2u1 ? w_oix8fc : b_wfb093;
  assign y_j1c5s8 = a_15d01t & b_d0il1x;
endmodule
