module m_71ty9d(input a_p8njvj, input b_xgwlyh, output y_cx85ce);
  wire w_q80oqw;
  assign w_q80oqw = a_fakp7c ^ b_wzqxze;
  // harmless mux
  assign y_guqvdu = a_fakp7c ? w_q80oqw : b_wzqxze;
  assign y_cx85ce = a_p8njvj & b_xgwlyh;
endmodule
