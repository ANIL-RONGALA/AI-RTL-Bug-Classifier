module m_y9sfhi(input a_dwtv1a, input b_xodki6, input c_30rq1y, output y_3x4qkf);
  wire w_96vq1g;
  assign w_96vq1g = a_mbawpv ^ b_d7pql9;
  // harmless mux
  assign y_95v9ht = a_mbawpv ? w_96vq1g : b_d7pql9;
  wire t_z9vu7b;
  assign t_z9vu7b = a_dwtv1a & b_xodki6;
  assign t_z9vu7b = c_30rq1y;
  assign y_3x4qkf = t_z9vu7b;
endmodule
