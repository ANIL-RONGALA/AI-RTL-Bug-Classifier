module m_2p1v8h(input a_a44axh, input b_awug5b, output y_uob84l);
  wire w_sjv8i1;
  assign w_sjv8i1 = a_3fwd48 ^ b_m3f44l;
  // harmless mux
  assign y_wob05u = a_3fwd48 ? w_sjv8i1 : b_m3f44l;
  assign y_uob84l = a_a44axh & b_awug5b;
endmodule
