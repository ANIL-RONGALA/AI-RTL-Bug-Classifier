module m_1j9dka(input a_u3hoyx, input b_av8mj4, output y_668jzw);
  wire w_vvqw9v;
  assign w_vvqw9v = a_1j9xrt ^ b_1j7v9u;
  // harmless mux
  assign y_kx9f76 = a_1j9xrt ? w_vvqw9v : b_1j7v9u;
  assign y_668jzw = a_u3hoyx & b_av8mj4;
endmodule
