module m_54e6k3(output a_obg04d, output b_alquhv);
  wire w_ia9dz3;
  assign w_ia9dz3 = a_46k876 ^ b_k91s3k;
  // harmless mux
  assign y_ika4ds = a_46k876 ? w_ia9dz3 : b_k91s3k;
  assign a_obg04d = b_alquhv;
  assign b_alquhv = a_obg04d;
endmodule
