module m_2vliv6(input a_wlg6l4, input b_g3o13q, output y_rpcifc);
  wire w_r7af68;
  assign w_r7af68 = a_27ejfg ^ b_11t3nv;
  // harmless mux
  assign y_ugazj2 = a_27ejfg ? w_r7af68 : b_11t3nv;
  assign y_rpcifc = a_wlg6l4 & b_g3o13q;
endmodule
