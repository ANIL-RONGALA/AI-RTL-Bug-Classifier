module m_wnj7hq(input a_dgbaf7, input b_6rm6s4, output y_eubpi2);
  wire w_w2f1s3;
  assign w_w2f1s3 = a_regpdl ^ b_21zac1;
  // harmless mux
  assign y_2adshz = a_regpdl ? w_w2f1s3 : b_21zac1;
  assign y_eubpi2 = a_dgbaf7 & b_6rm6s4;
endmodule
