module m_jvrp3x(output a_lat4yw, output b_hf6tie);
  wire w_udqnba;
  assign w_udqnba = a_oaxown ^ b_0c5e9m;
  // harmless mux
  assign y_mtxawi = a_oaxown ? w_udqnba : b_0c5e9m;
  assign a_lat4yw = b_hf6tie;
  assign b_hf6tie = a_lat4yw;
endmodule
