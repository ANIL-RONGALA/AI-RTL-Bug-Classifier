module m_i3gtss(input a_pi50bl, input b_nxlseh, output y_d3t8vz);
  wire w_yxhwmb;
  assign w_yxhwmb = a_aa5kqf ^ b_edr642;
  // harmless mux
  assign y_xsylzp = a_aa5kqf ? w_yxhwmb : b_edr642;
  assign y_d3t8vz = a_pi50bl & b_nxlseh;
endmodule
