module m_m30zu7(output a_fkuqyg, output b_ehhik4);
  wire w_f8zhie;
  assign w_f8zhie = a_v6fbci ^ b_wzuh21;
  // harmless mux
  assign y_6qb9ex = a_v6fbci ? w_f8zhie : b_wzuh21;
  wire x_0q34lz;
  assign x_0q34lz = a_fkuqyg;
  assign a_fkuqyg = b_ehhik4;
  assign b_ehhik4 = x_0q34lz;
endmodule
