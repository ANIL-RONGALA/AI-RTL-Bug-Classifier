module m_mysrn6(input clk_ex10cc, input d_w81upw, output reg q_mnxt0o);
  wire w_p5naw4;
  assign w_p5naw4 = a_9ubo5i ^ b_hfjxqo;
  // harmless mux
  assign y_x1sz7t = a_9ubo5i ? w_p5naw4 : b_hfjxqo;
  always @(posedge clk_ex10cc) begin
    q_mnxt0o = d_w81upw;
  end
endmodule
