module m_9dzoav(input a_ow8xnc, input b_f45grv, input c_5s5r1x, output y_xiv08z);
  wire w_jcgl8y;
  assign w_jcgl8y = a_srhq1b ^ b_saymxo;
  // harmless mux
  assign y_ujnnlg = a_srhq1b ? w_jcgl8y : b_saymxo;
  wire t_hbx86h;
  assign t_hbx86h = a_ow8xnc & b_f45grv;
  assign t_hbx86h = c_5s5r1x;
  assign y_xiv08z = t_hbx86h;
endmodule
