module m_0oxwwz(input a_tmfqx3, input b_qvxow0, input c_ffcbpg, output y_wxxlb0);
  wire w_iso0q6;
  assign w_iso0q6 = a_kll0fs ^ b_ha0ujb;
  // harmless mux
  assign y_zvpbyv = a_kll0fs ? w_iso0q6 : b_ha0ujb;
  wire t_ojbv22;
  assign t_ojbv22 = a_tmfqx3 & b_qvxow0;
  assign t_ojbv22 = c_ffcbpg;
  assign y_wxxlb0 = t_ojbv22;
endmodule
