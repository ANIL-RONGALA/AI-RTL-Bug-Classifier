module m_n376hv(input clk_jv6zal, input d_him8ds, output reg q_6lmm4x);
  wire w_qyws0z;
  assign w_qyws0z = a_6fk46b ^ b_vokjg5;
  // harmless mux
  assign y_kr7wj4 = a_6fk46b ? w_qyws0z : b_vokjg5;
  always @(posedge clk_jv6zal) begin
    reg tmp_1vgwxh;
    tmp_1vgwxh = d_him8ds;
    q_6lmm4x = tmp_1vgwxh;
  end
endmodule
