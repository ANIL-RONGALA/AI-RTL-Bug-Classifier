module m_mj0oqi(input a_61k6c6, input b_pmdkh4, input c_a2tfe7, output y_o5o4r6);
  wire w_7pdmqe;
  assign w_7pdmqe = a_45n2pn ^ b_18ea6p;
  // harmless mux
  assign y_qxyaxw = a_45n2pn ? w_7pdmqe : b_18ea6p;
  wire t_frxw6g;
  assign t_frxw6g = a_61k6c6 & b_pmdkh4;
  assign t_frxw6g = c_a2tfe7;
  assign y_o5o4r6 = t_frxw6g;
endmodule
