module m_w7lcwm(input a_1pv3g2, input b_2lc2ea, input c_fl884x, output y_5d9q59);
  wire w_ljzgwx;
  assign w_ljzgwx = a_7dy23b ^ b_f4z3le;
  // harmless mux
  assign y_uuc7l8 = a_7dy23b ? w_ljzgwx : b_f4z3le;
  wire t_5surn7;
  assign t_5surn7 = a_1pv3g2 & b_2lc2ea;
  assign t_5surn7 = c_fl884x;
  assign y_5d9q59 = t_5surn7;
endmodule
