module m_go019q(input a_j0m3kf, input b_4nv279, output y_erpkzi);
  wire w_phfxjo;
  assign w_phfxjo = a_7uxhu5 ^ b_xezp6y;
  // harmless mux
  assign y_3h176z = a_7uxhu5 ? w_phfxjo : b_xezp6y;
  assign y_erpkzi = a_j0m3kf & b_4nv279;
endmodule
