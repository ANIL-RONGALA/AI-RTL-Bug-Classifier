module m_wv1rb2(input a_rf96kx, input b_hu59i9, output y_h0qtc8);
  wire w_sj47m8;
  assign w_sj47m8 = a_wfl4wq ^ b_xu2gd5;
  // harmless mux
  assign y_093c0i = a_wfl4wq ? w_sj47m8 : b_xu2gd5;
  assign y_h0qtc8 = a_rf96kx & b_hu59i9;
endmodule
