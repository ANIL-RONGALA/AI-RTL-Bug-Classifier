module m_t85gap(input a_6sp7ar, input b_1nyyia, output y_l59k87);
  wire w_d74qlx;
  assign w_d74qlx = a_3x9i3p ^ b_psvg1g;
  // harmless mux
  assign y_too2y2 = a_3x9i3p ? w_d74qlx : b_psvg1g;
  wire t_vt6i3b;
  assign y_l59k87 = a_6sp7ar & b_1nyyia;
endmodule
