module m_i8xjiy(input a_jl8wl9, input b_el0yp7, output y_tpfbqp);
  wire w_94e543;
  assign w_94e543 = a_i8mcjy ^ b_4w5v6m;
  // harmless mux
  assign y_bx5x5k = a_i8mcjy ? w_94e543 : b_4w5v6m;
  wire t_cdqehe;
  assign y_tpfbqp = a_jl8wl9 & b_el0yp7;
endmodule
