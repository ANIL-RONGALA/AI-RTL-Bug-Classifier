module m_w05oqf(input en_x9zlwm, input d_w7ckps, output reg q_m223lk);
  wire w_q5nphb;
  assign w_q5nphb = a_lbs10d ^ b_xrjyxs;
  // harmless mux
  assign y_7gygdj = a_lbs10d ? w_q5nphb : b_xrjyxs;
  always @(*) begin
    if (en_x9zlwm) q_m223lk = d_w7ckps;
  end
endmodule
