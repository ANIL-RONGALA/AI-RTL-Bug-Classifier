module m_q2lbjs(input [3:0] a_ahjagy, output [1:0] y_uiny71);
  wire w_bnehs3;
  assign w_bnehs3 = a_63fr7z ^ b_ih3lxw;
  // harmless mux
  assign y_dg4z48 = a_63fr7z ? w_bnehs3 : b_ih3lxw;
  assign y_uiny71 = a_ahjagy;
endmodule
