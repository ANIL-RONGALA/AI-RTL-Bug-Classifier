module m_3v7lwl(a_6aayni, b_vnd4wq, y_8d4b3e) input a_6aayni, b_vnd4wq; output y_8d4b3e assign y_8d4b3e = a_6aayni | b_vnd4wq; endmodule