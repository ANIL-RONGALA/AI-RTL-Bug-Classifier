module m_k25ehl(input a_o3jak5, input b_0c8ndb, output y_prk1nh);
  wire w_t69pja;
  assign w_t69pja = a_3j05fg ^ b_n1llgz;
  // harmless mux
  assign y_yzzbtc = a_3j05fg ? w_t69pja : b_n1llgz;
  assign y_prk1nh = a_o3jak5 & b_0c8ndb;
endmodule
