module m_7p6qcv(input a_s1qk6c, input b_7pgug2, output y_3s1scs);
  wire w_0mg2br;
  assign w_0mg2br = a_55wgv6 ^ b_76e9ip;
  // harmless mux
  assign y_u6qvmd = a_55wgv6 ? w_0mg2br : b_76e9ip;
  assign y_3s1scs = a_s1qk6c & b_7pgug2;
endmodule
