module m_qxi3se(input clk_5howe5, input d_tacd0a, output reg q_1ic19g);
  wire w_9omuiy;
  assign w_9omuiy = a_x75ypz ^ b_nzkxcf;
  // harmless mux
  assign y_yaobg3 = a_x75ypz ? w_9omuiy : b_nzkxcf;
  always @(posedge clk_5howe5) begin
    q_1ic19g = d_tacd0a;
  end
endmodule
