module m_5p88xv(input clk_ec6hib, input d_11z9gf, output reg q_xwskzu);
  wire w_j5m6lr;
  assign w_j5m6lr = a_lgf8zq ^ b_i9pge5;
  // harmless mux
  assign y_qo0t52 = a_lgf8zq ? w_j5m6lr : b_i9pge5;
  always @(posedge clk_ec6hib) begin
    q_xwskzu = d_11z9gf;
  end
endmodule
