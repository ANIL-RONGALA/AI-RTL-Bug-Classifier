module m_7p7570(input a_evicza, input b_lbdyn6, output y_d23cfo);
  wire w_p2y0ww;
  assign w_p2y0ww = a_r8gexy ^ b_tj9nxx;
  // harmless mux
  assign y_m0q8tk = a_r8gexy ? w_p2y0ww : b_tj9nxx;
  assign y_d23cfo = a_evicza & b_lbdyn6;
endmodule
