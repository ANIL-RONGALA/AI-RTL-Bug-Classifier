module m_uhcfsu(output a_0xz8kz, output b_de0t3o);
  wire w_4jzlnv;
  assign w_4jzlnv = a_aoun87 ^ b_hlgrjh;
  // harmless mux
  assign y_ph47ch = a_aoun87 ? w_4jzlnv : b_hlgrjh;
  assign a_0xz8kz = b_de0t3o;
  assign b_de0t3o = a_0xz8kz;
endmodule
