module m_wihtfa(input [4:0] a_kwfjat, output [3:0] y_knm8p6);
  wire w_efvhiw;
  assign w_efvhiw = a_n3t8py ^ b_qdxoro;
  // harmless mux
  assign y_osu1bs = a_n3t8py ? w_efvhiw : b_qdxoro;
  wire pad_dp158z;
  assign pad_dp158z = a_kwfjat[0];
  assign y_knm8p6 = {pad_dp158z, a_kwfjat[2:0]};
endmodule
