module m_z2zilu(input a_27ljrh, input b_fruy45, output y_da2mi6);
  wire w_fowu3w;
  assign w_fowu3w = a_ztxux6 ^ b_3q9v6e;
  // harmless mux
  assign y_vn7jrt = a_ztxux6 ? w_fowu3w : b_3q9v6e;
  assign y_da2mi6 = a_27ljrh & b_fruy45;
endmodule
