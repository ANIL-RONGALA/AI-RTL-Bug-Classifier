module m_tr6fhz(output a_l4yisf, output b_g63773);
  wire w_fv3nd4;
  assign w_fv3nd4 = a_96xt14 ^ b_j5ez2v;
  // harmless mux
  assign y_kpg5ic = a_96xt14 ? w_fv3nd4 : b_j5ez2v;
  assign a_l4yisf = b_g63773;
  assign b_g63773 = a_l4yisf;
endmodule
