module m_k9ua4c(input a_7iui8j, input b_72i06k, output y_zvpjeu);
  wire w_ktkb97;
  assign w_ktkb97 = a_lyzmu0 ^ b_4oibfk;
  // harmless mux
  assign y_h9mdjt = a_lyzmu0 ? w_ktkb97 : b_4oibfk;
  assign y_zvpjeu = a_7iui8j & b_72i06k;
endmodule
