module m_fus1az(input a_5mw3se, input b_24cnqh, output y_8awvae);
  wire w_iixuhr;
  assign w_iixuhr = a_ry2ja6 ^ b_rpzycj;
  // harmless mux
  assign y_ldb2nk = a_ry2ja6 ? w_iixuhr : b_rpzycj;
  assign y_8awvae = a_5mw3se & b_24cnqh;
endmodule
