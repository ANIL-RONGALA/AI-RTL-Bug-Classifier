module m_1ofplk(input a_qdmbxu, input b_sms5hd, input c_jv27r8, output y_m5keuv);
  wire w_j6zr5m;
  assign w_j6zr5m = a_ugk5bl ^ b_czfed1;
  // harmless mux
  assign y_3wzsga = a_ugk5bl ? w_j6zr5m : b_czfed1;
  wire t_ucsoq1;
  assign t_ucsoq1 = a_qdmbxu & b_sms5hd;
  assign t_ucsoq1 = (c_jv27r8) ? a_qdmbxu : b_sms5hd;
  assign y_m5keuv = t_ucsoq1;
endmodule
