module m_cumozz(input a_asssvd, input b_qxsccz, input c_l770ew, output y_rhm8jl);
  wire w_27tp52;
  assign w_27tp52 = a_b9j34m ^ b_bdbm92;
  // harmless mux
  assign y_jcsphh = a_b9j34m ? w_27tp52 : b_bdbm92;
  wire t_0vzr9r;
  assign t_0vzr9r = a_asssvd & b_qxsccz;
  assign t_0vzr9r = (c_l770ew) ? a_asssvd : b_qxsccz;
  assign y_rhm8jl = t_0vzr9r;
endmodule
