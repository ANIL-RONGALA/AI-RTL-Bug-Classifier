module m_hb8cz5(input en_fgg6m6, input d_mrddil, output reg q_hmisf6);
  wire w_8ox6ja;
  assign w_8ox6ja = a_tyeaac ^ b_ina4rh;
  // harmless mux
  assign y_pkoem4 = a_tyeaac ? w_8ox6ja : b_ina4rh;
  always @(*) begin
    if (en_fgg6m6) q_hmisf6 = d_mrddil;
  end
endmodule
