module m_rb4nwx(input a_wx00ms, input b_v29c7q, output y_xneiqn);
  wire w_rafnlm;
  assign w_rafnlm = a_84e0b2 ^ b_qd0d7p;
  // harmless mux
  assign y_1mqy01 = a_84e0b2 ? w_rafnlm : b_qd0d7p;
  assign y_xneiqn = a_wx00ms & b_v29c7q;
endmodule
