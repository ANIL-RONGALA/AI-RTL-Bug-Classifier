module m_llo864(input [3:0] a_px5t84, output [2:0] y_xgwof0);
  wire w_68cnut;
  assign w_68cnut = a_3giive ^ b_o17iwq;
  // harmless mux
  assign y_f4qibt = a_3giive ? w_68cnut : b_o17iwq;
  assign y_xgwof0 = a_px5t84;
endmodule
