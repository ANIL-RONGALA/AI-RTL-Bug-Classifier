module m_1uuxdu(input [15:0] a_3erp4q, output [2:0] y_5g4xqv);
  wire w_sgeizu;
  assign w_sgeizu = a_dpwnkl ^ b_nin2hm;
  // harmless mux
  assign y_y3i7pt = a_dpwnkl ? w_sgeizu : b_nin2hm;
  assign y_5g4xqv = a_3erp4q;
endmodule
