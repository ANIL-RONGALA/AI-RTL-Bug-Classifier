module m_l3eszj(input a_po37gq, input b_fi4pm7, output y_pxospg);
  wire w_p0orqo;
  assign w_p0orqo = a_bhods3 ^ b_xfvgwl;
  // harmless mux
  assign y_ko0sge = a_bhods3 ? w_p0orqo : b_xfvgwl;
  assign y_pxospg = a_po37gq & b_fi4pm7;
endmodule
