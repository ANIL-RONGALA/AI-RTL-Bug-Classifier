module m_femflb(input a_jzgsv4, input b_ahr2rs, output y_k1mc8f);
  wire w_k5i9js;
  assign w_k5i9js = a_luwzm8 ^ b_j7sg23;
  // harmless mux
  assign y_8xzxiu = a_luwzm8 ? w_k5i9js : b_j7sg23;
  assign y_k1mc8f = a_jzgsv4 & b_ahr2rs;
endmodule
