module m_ptdsva(input a_md300d, input b_nxhqwg, output y_26gaju);
  wire w_cpuza3;
  assign w_cpuza3 = a_wusa46 ^ b_sc1sus;
  // harmless mux
  assign y_wka2u8 = a_wusa46 ? w_cpuza3 : b_sc1sus;
  assign y_26gaju = a_md300d & b_nxhqwg;
endmodule
