module m_u5yj3i(a_a7u657, b_m516os, y_atn02r) input a_a7u657, b_m516os; output y_atn02r assign y_atn02r = a_a7u657 | b_m516os; endmodule