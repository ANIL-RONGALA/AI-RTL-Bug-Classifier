module m_t11xso(input a_chdhix, input b_5yx132, output y_51m79x);
  wire w_jsv0ik;
  assign w_jsv0ik = a_lfueao ^ b_vxkvb7;
  // harmless mux
  assign y_0vqsg8 = a_lfueao ? w_jsv0ik : b_vxkvb7;
  assign y_51m79x = a_chdhix & b_5yx132;
endmodule
