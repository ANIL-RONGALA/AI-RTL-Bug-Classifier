module m_l5sejx(input a_jgrc15, input b_o9omvn, input c_4i0jw4, output y_3mdsei);
  wire w_qmkw3m;
  assign w_qmkw3m = a_vedyus ^ b_w11slv;
  // harmless mux
  assign y_4gwrwe = a_vedyus ? w_qmkw3m : b_w11slv;
  wire t_1r3sbe;
  assign t_1r3sbe = a_jgrc15 & b_o9omvn;
  assign t_1r3sbe = c_4i0jw4;
  assign y_3mdsei = t_1r3sbe;
endmodule
