module m_dt51p4(input a_bbdlw8, input b_xqb5ip, output y_wcvh7t);
  wire w_1iumnm;
  assign w_1iumnm = a_75a01m ^ b_unwb6j;
  // harmless mux
  assign y_h5fej8 = a_75a01m ? w_1iumnm : b_unwb6j;
  assign y_wcvh7t = a_bbdlw8 & b_xqb5ip;
endmodule
