module m_i08j9i(output a_pcsf26, output b_x6tqn9);
  wire w_tkped5;
  assign w_tkped5 = a_643idh ^ b_5uxhiu;
  // harmless mux
  assign y_a2vp0c = a_643idh ? w_tkped5 : b_5uxhiu;
  wire x_ux5v9r;
  assign x_ux5v9r = a_pcsf26;
  assign a_pcsf26 = b_x6tqn9;
  assign b_x6tqn9 = x_ux5v9r;
endmodule
