module m_93b7ie(input a_ldc4jz, input b_371hh7, output y_73klez);
  wire w_vly7b6;
  assign w_vly7b6 = a_s74f4g ^ b_3ptukt;
  // harmless mux
  assign y_gmv3qs = a_s74f4g ? w_vly7b6 : b_3ptukt;
  assign y_73klez = a_ldc4jz & b_371hh7;
endmodule
