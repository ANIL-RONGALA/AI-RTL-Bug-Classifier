module m_5zx7fs(output a_ookaqx, output b_b84pbr);
  wire w_vx9k3p;
  assign w_vx9k3p = a_dq2i7p ^ b_a0aro1;
  // harmless mux
  assign y_14vya7 = a_dq2i7p ? w_vx9k3p : b_a0aro1;
  wire x_s3gvk9;
  assign x_s3gvk9 = a_ookaqx;
  assign a_ookaqx = b_b84pbr;
  assign b_b84pbr = x_s3gvk9;
endmodule
