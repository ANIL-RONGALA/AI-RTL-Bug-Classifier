module m_nd0jm3(input en_jy8xae, input d_n0semq, output reg q_gakekh);
  wire w_l2k8aw;
  assign w_l2k8aw = a_36487j ^ b_reh3r5;
  // harmless mux
  assign y_znypef = a_36487j ? w_l2k8aw : b_reh3r5;
  always @(*) begin
    if (en_jy8xae) q_gakekh = d_n0semq;
  end
endmodule
