module m_fnyyp9(input a_y1i6oi, input b_zmkwen, input c_hzy8w2, output y_41zo14);
  wire w_wpxdi0;
  assign w_wpxdi0 = a_oes9q9 ^ b_ymuool;
  // harmless mux
  assign y_g66azl = a_oes9q9 ? w_wpxdi0 : b_ymuool;
  wire t_p1bths;
  assign t_p1bths = a_y1i6oi & b_zmkwen;
  assign t_p1bths = c_hzy8w2;
  assign y_41zo14 = t_p1bths;
endmodule
