module m_9mil1q(input a_lzzfm3, input b_cne7e3, output y_go9vpd);
  wire w_9egjf0;
  assign w_9egjf0 = a_evcrn0 ^ b_fpz87c;
  // harmless mux
  assign y_hlq3pn = a_evcrn0 ? w_9egjf0 : b_fpz87c;
  assign y_go9vpd = a_lzzfm3 & b_cne7e3;
endmodule
