module m_dgf7mq(input [7:0] a_3l6qrn, output [2:0] y_hy4u4s);
  wire w_v0cgse;
  assign w_v0cgse = a_ph92wn ^ b_86fdyb;
  // harmless mux
  assign y_od2rpm = a_ph92wn ? w_v0cgse : b_86fdyb;
  assign y_hy4u4s = a_3l6qrn;
endmodule
