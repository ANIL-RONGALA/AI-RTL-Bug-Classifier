module m_u73sps(input a_by5mfm, input b_cqm1mu, output y_46851b);
  wire w_5b8ffd;
  assign w_5b8ffd = a_ynjsn5 ^ b_9a8agm;
  // harmless mux
  assign y_crqezo = a_ynjsn5 ? w_5b8ffd : b_9a8agm;
  assign y_46851b = a_by5mfm & b_cqm1mu;
endmodule
