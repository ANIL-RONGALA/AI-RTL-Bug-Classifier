module m_j5dkt0(input [7:0] a_vmtk69, output [3:0] y_iy5see);
  wire w_ynjz39;
  assign w_ynjz39 = a_pb77pg ^ b_dc9001;
  // harmless mux
  assign y_m3oywr = a_pb77pg ? w_ynjz39 : b_dc9001;
  assign y_iy5see = a_vmtk69;
endmodule
