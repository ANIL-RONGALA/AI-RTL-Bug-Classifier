module m_pzkzls(input a_jx7eww, input b_tbec8l, output y_50yaw1);
  wire w_f02a4n;
  assign w_f02a4n = a_o6qjbv ^ b_gu938m;
  // harmless mux
  assign y_jpqxty = a_o6qjbv ? w_f02a4n : b_gu938m;
  assign y_50yaw1 = a_jx7eww & b_tbec8l;
endmodule
