module m_yn5bqw(input a_rsjdsq, input b_czigg5, output y_1xm1vz);
  wire w_vm1uxa;
  assign w_vm1uxa = a_gyhtdw ^ b_nhqxg2;
  // harmless mux
  assign y_rp5oow = a_gyhtdw ? w_vm1uxa : b_nhqxg2;
  wire t_he5b8m;
  assign t_he5b8m = a_rsjdsq | b_czigg5;
  assign y_1xm1vz = a_rsjdsq & b_czigg5;
endmodule
