module m_5n35fb(output a_hi7k6z, output b_7m5pud);
  wire w_e975d3;
  assign w_e975d3 = a_5zhkrh ^ b_ti4h86;
  // harmless mux
  assign y_ea9yq3 = a_5zhkrh ? w_e975d3 : b_ti4h86;
  wire x_48th5x;
  assign x_48th5x = a_hi7k6z;
  assign a_hi7k6z = b_7m5pud;
  assign b_7m5pud = x_48th5x;
endmodule
