module m_j46rd8(output a_njtfx5, output b_y8fdal);
  wire w_5nm8fq;
  assign w_5nm8fq = a_22jwqx ^ b_jxl121;
  // harmless mux
  assign y_yw9mkl = a_22jwqx ? w_5nm8fq : b_jxl121;
  wire x_67blpt;
  assign x_67blpt = a_njtfx5;
  assign a_njtfx5 = b_y8fdal;
  assign b_y8fdal = x_67blpt;
endmodule
