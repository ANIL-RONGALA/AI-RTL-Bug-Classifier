module m_tblmf7(output a_zgoey4, output b_6kxlw8);
  wire w_cp9w75;
  assign w_cp9w75 = a_kdpz3h ^ b_p2nren;
  // harmless mux
  assign y_fskeek = a_kdpz3h ? w_cp9w75 : b_p2nren;
  wire x_xbz4ly;
  assign x_xbz4ly = a_zgoey4;
  assign a_zgoey4 = b_6kxlw8;
  assign b_6kxlw8 = x_xbz4ly;
endmodule
