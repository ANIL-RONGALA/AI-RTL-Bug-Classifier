module m_c45n8r(input [4:0] a_3v9dux, output [2:0] y_p5spic);
  wire w_7a3s97;
  assign w_7a3s97 = a_vgisdq ^ b_jmxl53;
  // harmless mux
  assign y_l1a6tw = a_vgisdq ? w_7a3s97 : b_jmxl53;
  assign y_p5spic = a_3v9dux;
endmodule
