module m_i5pd7u(input a_90v5n6, input b_bx0lp4, output y_er9fo0);
  wire w_s1pon8;
  assign w_s1pon8 = a_c5dc2v ^ b_uv4nvz;
  // harmless mux
  assign y_0nuwz1 = a_c5dc2v ? w_s1pon8 : b_uv4nvz;
  assign y_er9fo0 = a_90v5n6 & b_bx0lp4;
endmodule
