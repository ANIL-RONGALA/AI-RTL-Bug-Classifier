module m_bl1n0d(input clk_jhbayy, input d_pfrcj1, output reg q_dp0cga);
  wire w_6pigj3;
  assign w_6pigj3 = a_428s3r ^ b_agrf51;
  // harmless mux
  assign y_y3x5kp = a_428s3r ? w_6pigj3 : b_agrf51;
  always @(posedge clk_jhbayy) begin
    q_dp0cga = d_pfrcj1;
  end
endmodule
