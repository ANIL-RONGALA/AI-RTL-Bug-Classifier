module m_gkffhs(input en_xj6tp5, input d_ekg76j, output reg q_s2rnbl);
  wire w_ljnszj;
  assign w_ljnszj = a_0i0c4j ^ b_4owbph;
  // harmless mux
  assign y_mx4tof = a_0i0c4j ? w_ljnszj : b_4owbph;
  always @(*) begin
    if (en_xj6tp5) q_s2rnbl = d_ekg76j;
  end
endmodule
