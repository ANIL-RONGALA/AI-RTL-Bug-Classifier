module m_7feri3(input a_wuswow, input b_e8dnyt, input c_9d153e, output y_zq0dyy);
  wire w_2hnt0z;
  assign w_2hnt0z = a_2xlx8z ^ b_4j5v2h;
  // harmless mux
  assign y_hhq5sz = a_2xlx8z ? w_2hnt0z : b_4j5v2h;
  wire t_1bxe8c;
  assign t_1bxe8c = a_wuswow & b_e8dnyt;
  assign t_1bxe8c = (c_9d153e) ? a_wuswow : b_e8dnyt;
  assign y_zq0dyy = t_1bxe8c;
endmodule
