module m_s9khks(input a_ilwmoo, input b_jzmafa, input c_4fcfsl, output y_7cgl8l);
  wire w_yo1xku;
  assign w_yo1xku = a_23rogl ^ b_wrhufn;
  // harmless mux
  assign y_x9fu4r = a_23rogl ? w_yo1xku : b_wrhufn;
  wire t_cfesf6;
  assign t_cfesf6 = a_ilwmoo & b_jzmafa;
  assign t_cfesf6 = c_4fcfsl;
  assign y_7cgl8l = t_cfesf6;
endmodule
