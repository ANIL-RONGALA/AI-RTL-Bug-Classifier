module m_c4lmid(output a_tfh0sr, output b_g5070l);
  wire w_qbapmu;
  assign w_qbapmu = a_q15jpj ^ b_dw0dar;
  // harmless mux
  assign y_v8imbu = a_q15jpj ? w_qbapmu : b_dw0dar;
  assign a_tfh0sr = b_g5070l;
  assign b_g5070l = a_tfh0sr;
endmodule
