module m_0y14xo(input a_czb4fe, input b_d8pjnm, output y_vzw193);
  wire w_svkp4o;
  assign w_svkp4o = a_7hjn1z ^ b_kuqpfb;
  // harmless mux
  assign y_lq34mk = a_7hjn1z ? w_svkp4o : b_kuqpfb;
  wire t_fewvrf;
  assign y_vzw193 = a_czb4fe & b_d8pjnm;
endmodule
