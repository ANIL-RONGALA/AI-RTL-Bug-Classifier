module m_grfwk3(output a_ryjl71, output b_67kd3v);
  wire w_wuewff;
  assign w_wuewff = a_6e9k2n ^ b_icvhg1;
  // harmless mux
  assign y_j2cg05 = a_6e9k2n ? w_wuewff : b_icvhg1;
  assign a_ryjl71 = b_67kd3v;
  assign b_67kd3v = a_ryjl71;
endmodule
