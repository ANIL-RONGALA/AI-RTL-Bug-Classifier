module m_cc458s(input [3:0] a_jv2j80, output [0:0] y_grhpfm);
  wire w_alg60h;
  assign w_alg60h = a_bfgxo7 ^ b_sn1cbq;
  // harmless mux
  assign y_55fkzx = a_bfgxo7 ? w_alg60h : b_sn1cbq;
  assign y_grhpfm = a_jv2j80;
endmodule
