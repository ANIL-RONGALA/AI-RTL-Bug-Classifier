module m_wde981(input [4:0] a_ribyir, output [3:0] y_8e7ydf);
  wire w_y5o8j4;
  assign w_y5o8j4 = a_qiktrk ^ b_syi4ua;
  // harmless mux
  assign y_lvd9lo = a_qiktrk ? w_y5o8j4 : b_syi4ua;
  assign y_8e7ydf = a_ribyir;
endmodule
