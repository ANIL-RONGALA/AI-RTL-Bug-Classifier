module m_t8anon(input a_vew0yb, input b_uubkap, output y_8u8ay8);
  wire w_mx6759;
  assign w_mx6759 = a_ohbeu6 ^ b_kznqi0;
  // harmless mux
  assign y_f42d57 = a_ohbeu6 ? w_mx6759 : b_kznqi0;
  wire t_ntprw8;
  assign y_8u8ay8 = a_vew0yb & b_uubkap;
endmodule
