module m_58qwtk(input a_s1p5yv, input b_xm47um, output y_3ew1b4);
  wire w_fam2d8;
  assign w_fam2d8 = a_7ycwvp ^ b_13f8fd;
  // harmless mux
  assign y_bo1fis = a_7ycwvp ? w_fam2d8 : b_13f8fd;
  assign y_3ew1b4 = a_s1p5yv & b_xm47um;
endmodule
