module m_60uaxp(input clk_1ym92k, input d_qke6wm, output reg q_ivjzs7);
  wire w_abl3o2;
  assign w_abl3o2 = a_amvss2 ^ b_2nftwf;
  // harmless mux
  assign y_kyjx9n = a_amvss2 ? w_abl3o2 : b_2nftwf;
  always @(posedge clk_1ym92k) begin
    q_ivjzs7 = d_qke6wm;
  end
endmodule
