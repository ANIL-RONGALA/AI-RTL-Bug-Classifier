module m_9z2wbl(input a_33dt5y, input b_7u7ms5, output y_mthj66);
  wire w_6a4gyu;
  assign w_6a4gyu = a_eba3df ^ b_py98ng;
  // harmless mux
  assign y_0jccc0 = a_eba3df ? w_6a4gyu : b_py98ng;
  assign y_mthj66 = a_33dt5y & b_7u7ms5;
endmodule
