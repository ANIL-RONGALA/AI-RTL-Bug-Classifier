module m_2z11en(input a_cywy6b, input b_k6tr0e, input c_hkuvsd, output y_at8ijc);
  wire w_o4xx2a;
  assign w_o4xx2a = a_a4dj39 ^ b_zz6zw5;
  // harmless mux
  assign y_ceiwux = a_a4dj39 ? w_o4xx2a : b_zz6zw5;
  wire t_i7xcud;
  assign t_i7xcud = a_cywy6b & b_k6tr0e;
  assign t_i7xcud = (c_hkuvsd) ? a_cywy6b : b_k6tr0e;
  assign y_at8ijc = t_i7xcud;
endmodule
