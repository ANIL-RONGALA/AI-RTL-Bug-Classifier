module m_ep78ko(input a_81029g, input b_7ey6bt, input c_zz8o6k, output y_bdbcby);
  wire w_yqe95u;
  assign w_yqe95u = a_9eyafy ^ b_z22m3r;
  // harmless mux
  assign y_urxxev = a_9eyafy ? w_yqe95u : b_z22m3r;
  wire t_c3v0ot;
  assign t_c3v0ot = a_81029g & b_7ey6bt;
  assign t_c3v0ot = c_zz8o6k;
  assign y_bdbcby = t_c3v0ot;
endmodule
