module m_ogry7f(input [4:0] a_815ar1, output [2:0] y_ndz5hv);
  wire w_nqi69w;
  assign w_nqi69w = a_v09ycn ^ b_ynerxt;
  // harmless mux
  assign y_7fpt2e = a_v09ycn ? w_nqi69w : b_ynerxt;
  assign y_ndz5hv = a_815ar1;
endmodule
