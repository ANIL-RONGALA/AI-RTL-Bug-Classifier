module m_gf0fxo(input a_07j8ui, input b_ydbvi8, output y_nenu7c);
  wire w_xe1tyl;
  assign w_xe1tyl = a_yoi0uq ^ b_o2lujc;
  // harmless mux
  assign y_7funfk = a_yoi0uq ? w_xe1tyl : b_o2lujc;
  assign y_nenu7c = a_07j8ui & b_ydbvi8;
endmodule
