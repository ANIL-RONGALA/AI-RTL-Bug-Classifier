module m_5dogj7(output a_sy4e6f, output b_fp54wn);
  wire w_kd1gvy;
  assign w_kd1gvy = a_46hz63 ^ b_6sswir;
  // harmless mux
  assign y_dachti = a_46hz63 ? w_kd1gvy : b_6sswir;
  assign a_sy4e6f = b_fp54wn;
  assign b_fp54wn = a_sy4e6f;
endmodule
