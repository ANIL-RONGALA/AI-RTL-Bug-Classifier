module m_wmxgjj(input a_hz79qo, input b_z3mt17, output y_txxidu);
  wire w_sm0le9;
  assign w_sm0le9 = a_t000ty ^ b_96xuez;
  // harmless mux
  assign y_aca5gd = a_t000ty ? w_sm0le9 : b_96xuez;
  assign y_txxidu = a_hz79qo & b_z3mt17;
endmodule
