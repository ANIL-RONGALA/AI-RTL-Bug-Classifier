module m_0w66ab(input a_qnrge6, input b_q0nmxi, input c_2azlzg, output y_3p5asn);
  wire w_x804tt;
  assign w_x804tt = a_n8siyt ^ b_4ppniy;
  // harmless mux
  assign y_p7je3r = a_n8siyt ? w_x804tt : b_4ppniy;
  wire t_cvyln0;
  assign t_cvyln0 = a_qnrge6 & b_q0nmxi;
  assign t_cvyln0 = (c_2azlzg) ? a_qnrge6 : b_q0nmxi;
  assign y_3p5asn = t_cvyln0;
endmodule
