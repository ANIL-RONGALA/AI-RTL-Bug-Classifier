module m_sbtzre(input a_r1bezc, input b_c47xlw, output y_l2zplx);
  wire w_ar1wl9;
  assign w_ar1wl9 = a_wk2ere ^ b_b5x3gt;
  // harmless mux
  assign y_txmf70 = a_wk2ere ? w_ar1wl9 : b_b5x3gt;
  assign y_l2zplx = a_r1bezc & b_c47xlw;
endmodule
