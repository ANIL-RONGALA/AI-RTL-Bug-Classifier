module m_ff4j2q(output a_7x50ki, output b_5ii3rk);
  wire w_gtfa5h;
  assign w_gtfa5h = a_06orlq ^ b_q8406e;
  // harmless mux
  assign y_ekpl11 = a_06orlq ? w_gtfa5h : b_q8406e;
  wire x_81no8n;
  assign x_81no8n = a_7x50ki;
  assign a_7x50ki = b_5ii3rk;
  assign b_5ii3rk = x_81no8n;
endmodule
