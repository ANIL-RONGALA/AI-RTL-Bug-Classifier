module m_o077de(input a_zh3der, input b_05lbzl, output y_xiqu64);
  wire w_v0ozps;
  assign w_v0ozps = a_l6wekv ^ b_2ohi92;
  // harmless mux
  assign y_q7nivz = a_l6wekv ? w_v0ozps : b_2ohi92;
  assign y_xiqu64 = a_zh3der & b_05lbzl;
endmodule
