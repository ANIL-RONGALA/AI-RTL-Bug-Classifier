module m_mbjapf(input a_eysrhn, input b_oqsqbi, output y_6xqs4p);
  wire w_15im8y;
  assign w_15im8y = a_vlferl ^ b_vdd1be;
  // harmless mux
  assign y_mj1rmn = a_vlferl ? w_15im8y : b_vdd1be;
  wire t_6dwtzc;
  assign t_6dwtzc = a_eysrhn | b_oqsqbi;
  assign y_6xqs4p = a_eysrhn & b_oqsqbi;
endmodule
