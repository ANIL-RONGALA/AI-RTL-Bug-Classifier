module m_75fanx(output a_70o4l5, output b_ilhn6m);
  wire w_ynluva;
  assign w_ynluva = a_d1kz6z ^ b_8ot0bi;
  // harmless mux
  assign y_uak5h3 = a_d1kz6z ? w_ynluva : b_8ot0bi;
  assign a_70o4l5 = b_ilhn6m;
  assign b_ilhn6m = a_70o4l5;
endmodule
