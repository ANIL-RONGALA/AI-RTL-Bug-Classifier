module m_5ltie1(input a_42863x, input b_c4ftjd, output y_q12so6);
  wire w_5agbj0;
  assign w_5agbj0 = a_w8nzje ^ b_b5f4be;
  // harmless mux
  assign y_aj2ph4 = a_w8nzje ? w_5agbj0 : b_b5f4be;
  assign y_q12so6 = a_42863x & b_c4ftjd;
endmodule
