module m_3kzjgo(input [15:0] a_45xjus, output [1:0] y_ft0kl9);
  wire w_ad7z53;
  assign w_ad7z53 = a_0zkuie ^ b_1o22pg;
  // harmless mux
  assign y_3xvwnz = a_0zkuie ? w_ad7z53 : b_1o22pg;
  wire pad_h7s2dx;
  assign pad_h7s2dx = a_45xjus[0];
  assign y_ft0kl9 = {pad_h7s2dx, a_45xjus[0:0]};
endmodule
