module m_ooycr6(input a_ghgjzp, input b_eylwmi, output y_4jbmwx);
  wire w_puwlen;
  assign w_puwlen = a_t9pd97 ^ b_zqnpla;
  // harmless mux
  assign y_b0yumn = a_t9pd97 ? w_puwlen : b_zqnpla;
  assign y_4jbmwx = a_ghgjzp & b_eylwmi;
endmodule
