module m_9rlegt(input a_stymj4, input b_dmbyq3, input c_rzskp9, output y_89zh91);
  wire w_d8pm8s;
  assign w_d8pm8s = a_bizh86 ^ b_r1ph9f;
  // harmless mux
  assign y_wrbf2r = a_bizh86 ? w_d8pm8s : b_r1ph9f;
  wire t_eud92h;
  assign t_eud92h = a_stymj4 & b_dmbyq3;
  assign t_eud92h = c_rzskp9;
  assign y_89zh91 = t_eud92h;
endmodule
