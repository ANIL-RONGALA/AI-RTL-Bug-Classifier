module m_z7vg6d(input a_kom12a, input b_ajstyc, input c_7bmnk6, output y_j7762l);
  wire w_n5mq0r;
  assign w_n5mq0r = a_jforkr ^ b_31m1r5;
  // harmless mux
  assign y_7ykawv = a_jforkr ? w_n5mq0r : b_31m1r5;
  wire t_6uesc7;
  assign t_6uesc7 = a_kom12a & b_ajstyc;
  assign t_6uesc7 = (c_7bmnk6) ? a_kom12a : b_ajstyc;
  assign y_j7762l = t_6uesc7;
endmodule
