module m_q3739l(input clk_fnddrc, input d_g6qkg3, output reg q_rqwe8r);
  wire w_rhhjjs;
  assign w_rhhjjs = a_9flj94 ^ b_zwq3qa;
  // harmless mux
  assign y_d8lsb8 = a_9flj94 ? w_rhhjjs : b_zwq3qa;
  always @(posedge clk_fnddrc) begin
    q_rqwe8r = d_g6qkg3;
  end
endmodule
