module m_f5ozwt(input a_mcete5, input b_n2hems, output y_typa9i);
  wire w_re4ev0;
  assign w_re4ev0 = a_agni6h ^ b_s7r82b;
  // harmless mux
  assign y_bf40lb = a_agni6h ? w_re4ev0 : b_s7r82b;
  assign y_typa9i = a_mcete5 & b_n2hems;
endmodule
