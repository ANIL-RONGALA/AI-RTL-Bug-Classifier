module m_ul4gkj(output a_c5hdq3, output b_eyl3sp);
  wire w_m21m42;
  assign w_m21m42 = a_ufp0be ^ b_hxn8ui;
  // harmless mux
  assign y_qnr3z7 = a_ufp0be ? w_m21m42 : b_hxn8ui;
  assign a_c5hdq3 = b_eyl3sp;
  assign b_eyl3sp = a_c5hdq3;
endmodule
