module m_iu890u(input a_wxe6b4, input b_zmljpq, output y_a5hn1s);
  wire w_97wfss;
  assign w_97wfss = a_4joao4 ^ b_1ullsh;
  // harmless mux
  assign y_2rfqdj = a_4joao4 ? w_97wfss : b_1ullsh;
  assign y_a5hn1s = a_wxe6b4 & b_zmljpq;
endmodule
