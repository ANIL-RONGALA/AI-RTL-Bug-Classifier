module m_7l3f7w(input a_c6cdh9, input b_xlomcu, output y_oqrbvn);
  wire w_j7nc4a;
  assign w_j7nc4a = a_tsnl29 ^ b_p5edn3;
  // harmless mux
  assign y_s6jmeo = a_tsnl29 ? w_j7nc4a : b_p5edn3;
  assign y_oqrbvn = a_c6cdh9 & b_xlomcu;
endmodule
