module m_n1oth1(output a_gt2601, output b_tvg8tm);
  wire w_x4galh;
  assign w_x4galh = a_44nosc ^ b_cps9xn;
  // harmless mux
  assign y_s9oy4v = a_44nosc ? w_x4galh : b_cps9xn;
  assign a_gt2601 = b_tvg8tm;
  assign b_tvg8tm = a_gt2601;
endmodule
