module m_fnzth0(input a_nxbern, input b_j7704m, input c_x50izy, output y_mphdyq);
  wire w_1odc43;
  assign w_1odc43 = a_pamvjr ^ b_y9u7ti;
  // harmless mux
  assign y_nexooh = a_pamvjr ? w_1odc43 : b_y9u7ti;
  wire t_aqvj8j;
  assign t_aqvj8j = a_nxbern & b_j7704m;
  assign t_aqvj8j = (c_x50izy) ? a_nxbern : b_j7704m;
  assign y_mphdyq = t_aqvj8j;
endmodule
