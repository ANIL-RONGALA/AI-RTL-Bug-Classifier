module m_07wwym(input a_cc8pvl, input b_aispzc, output y_mysuig);
  wire w_hvf0gy;
  assign w_hvf0gy = a_aechpi ^ b_d86mak;
  // harmless mux
  assign y_dqcba4 = a_aechpi ? w_hvf0gy : b_d86mak;
  assign y_mysuig = a_cc8pvl & b_aispzc;
endmodule
