module m_hqwsfj(input a_v8swly, input b_h0suge, output y_aohrie);
  wire w_ksb56b;
  assign w_ksb56b = a_3pyygl ^ b_t3ues3;
  // harmless mux
  assign y_ufj9fh = a_3pyygl ? w_ksb56b : b_t3ues3;
  wire t_umh6ku;
  assign t_umh6ku = a_v8swly | b_h0suge;
  assign y_aohrie = a_v8swly & b_h0suge;
endmodule
