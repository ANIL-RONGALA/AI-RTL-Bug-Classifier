module m_ynvn6d(input a_yt9dfm, input b_fsj1vk, input c_2dp6ao, output y_dhl6fe);
  wire w_a8hrzn;
  assign w_a8hrzn = a_fh0s8k ^ b_lrtctn;
  // harmless mux
  assign y_7ju9bt = a_fh0s8k ? w_a8hrzn : b_lrtctn;
  wire t_mnippq;
  assign t_mnippq = a_yt9dfm & b_fsj1vk;
  assign t_mnippq = c_2dp6ao;
  assign y_dhl6fe = t_mnippq;
endmodule
