module m_abfreo(input a_q5gw3s, input b_25i6z2, output y_mtbv5f);
  wire w_g96aw8;
  assign w_g96aw8 = a_tjhj8p ^ b_hmuao3;
  // harmless mux
  assign y_tgrlfb = a_tjhj8p ? w_g96aw8 : b_hmuao3;
  assign y_mtbv5f = a_q5gw3s & b_25i6z2;
endmodule
