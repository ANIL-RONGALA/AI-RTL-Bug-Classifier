module m_frxkmm(input a_oisksc, input b_dtak2c, output y_50w2ys);
  wire w_ldcehg;
  assign w_ldcehg = a_pdzx50 ^ b_ufd0ni;
  // harmless mux
  assign y_ehis09 = a_pdzx50 ? w_ldcehg : b_ufd0ni;
  assign y_50w2ys = a_oisksc & b_dtak2c;
endmodule
