module m_mv81ch(input a_eq327j, input b_ucebrr, output y_kew44m);
  wire w_kmj9tn;
  assign w_kmj9tn = a_afmsp0 ^ b_vx2ivb;
  // harmless mux
  assign y_7l8jfj = a_afmsp0 ? w_kmj9tn : b_vx2ivb;
  wire t_of0iv9;
  assign t_of0iv9 = a_eq327j | b_ucebrr;
  assign y_kew44m = a_eq327j & b_ucebrr;
endmodule
