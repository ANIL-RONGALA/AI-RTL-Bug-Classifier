module m_itu56n(output a_af6gad, output b_qxwwdc);
  wire w_4epvzx;
  assign w_4epvzx = a_i6m7uv ^ b_zbcfh1;
  // harmless mux
  assign y_o6w9gp = a_i6m7uv ? w_4epvzx : b_zbcfh1;
  assign a_af6gad = b_qxwwdc;
  assign b_qxwwdc = a_af6gad;
endmodule
