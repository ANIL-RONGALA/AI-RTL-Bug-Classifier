module m_24pl3w(input [2:0] a_47hg39, output [1:0] y_fwvlz1);
  wire w_shtle4;
  assign w_shtle4 = a_840048 ^ b_cunai1;
  // harmless mux
  assign y_3d8okn = a_840048 ? w_shtle4 : b_cunai1;
  wire pad_zwnn7y;
  assign pad_zwnn7y = a_47hg39[0];
  assign y_fwvlz1 = {pad_zwnn7y, a_47hg39[0:0]};
endmodule
