module m_9acq9z(input a_mnqnin, input b_gkr9fu, output y_8183ei);
  wire w_o0lml1;
  assign w_o0lml1 = a_cjo9sb ^ b_qukzqx;
  // harmless mux
  assign y_wxyl8c = a_cjo9sb ? w_o0lml1 : b_qukzqx;
  assign y_8183ei = a_mnqnin & b_gkr9fu;
endmodule
