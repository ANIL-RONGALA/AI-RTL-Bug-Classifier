module m_v6p2ry(input a_4qqzhy, input b_4o6i5i, output y_210y0k);
  wire w_fu4j5p;
  assign w_fu4j5p = a_rfzueh ^ b_ef97ll;
  // harmless mux
  assign y_gocmut = a_rfzueh ? w_fu4j5p : b_ef97ll;
  wire t_1muf2b;
  assign y_210y0k = a_4qqzhy & b_4o6i5i;
endmodule
