module m_ha7ted(input a_67asoz, input b_lp5zjt, output y_927s2c);
  wire w_5n4kan;
  assign w_5n4kan = a_99k1jd ^ b_ruqou5;
  // harmless mux
  assign y_ugxc3q = a_99k1jd ? w_5n4kan : b_ruqou5;
  assign y_927s2c = a_67asoz & b_lp5zjt;
endmodule
