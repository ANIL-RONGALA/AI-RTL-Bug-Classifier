module m_dpyz6u(input a_a1p96f, input b_ogaasj, output y_iceis1);
  wire w_3u4y0g;
  assign w_3u4y0g = a_4k3k4f ^ b_p8pmj8;
  // harmless mux
  assign y_44kwnp = a_4k3k4f ? w_3u4y0g : b_p8pmj8;
  assign y_iceis1 = a_a1p96f & b_ogaasj;
endmodule
