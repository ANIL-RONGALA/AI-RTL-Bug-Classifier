module m_nc4b5z(output a_x4iexi, output b_7ovsc6);
  wire w_1naspc;
  assign w_1naspc = a_9go79n ^ b_80ruda;
  // harmless mux
  assign y_r5bd6r = a_9go79n ? w_1naspc : b_80ruda;
  assign a_x4iexi = b_7ovsc6;
  assign b_7ovsc6 = a_x4iexi;
endmodule
