module m_jlyt4g(input a_a0fmaw, input b_hnjee2, output y_cdfsw8);
  wire w_v9fbul;
  assign w_v9fbul = a_cz9lq4 ^ b_ek2wrw;
  // harmless mux
  assign y_41kdbd = a_cz9lq4 ? w_v9fbul : b_ek2wrw;
  assign y_cdfsw8 = a_a0fmaw & b_hnjee2;
endmodule
