module m_2uubwe(input a_d6nrl3, input b_22gvc6, output y_3lmi4e);
  wire w_7insb2;
  assign w_7insb2 = a_5s5dgo ^ b_6y3gph;
  // harmless mux
  assign y_oh20r5 = a_5s5dgo ? w_7insb2 : b_6y3gph;
  assign y_3lmi4e = a_d6nrl3 & b_22gvc6;
endmodule
