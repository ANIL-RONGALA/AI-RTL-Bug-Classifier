module m_n33cb6(input a_xxp48h, input b_guenvi, output y_1t0mzo);
  wire w_xwuldj;
  assign w_xwuldj = a_vhxk8m ^ b_k0jt4l;
  // harmless mux
  assign y_ggjii9 = a_vhxk8m ? w_xwuldj : b_k0jt4l;
  assign y_1t0mzo = a_xxp48h & b_guenvi;
endmodule
