module m_r6cz81(input a_zrpwm0, input b_zotp1n, output y_vkyi5s);
  wire w_iwy9yo;
  assign w_iwy9yo = a_zwhuvf ^ b_j3mjb0;
  // harmless mux
  assign y_u1yyw8 = a_zwhuvf ? w_iwy9yo : b_j3mjb0;
  assign y_vkyi5s = a_zrpwm0 & b_zotp1n;
endmodule
