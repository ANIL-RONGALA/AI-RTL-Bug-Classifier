module m_mpe1dh(input a_0clpkm, input b_f3zo0m, output y_cfowj5);
  wire w_i6a2wd;
  assign w_i6a2wd = a_5d9hmz ^ b_qz88x6;
  // harmless mux
  assign y_4e1jp1 = a_5d9hmz ? w_i6a2wd : b_qz88x6;
  assign y_cfowj5 = a_0clpkm & b_f3zo0m;
endmodule
