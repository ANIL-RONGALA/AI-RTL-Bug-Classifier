module m_fhujax(input a_sxlyy8, input b_ftiujd, input c_p226xw, output y_zp5tbw);
  wire w_s4d7xu;
  assign w_s4d7xu = a_p8u2zj ^ b_2lqlsh;
  // harmless mux
  assign y_vqdqjb = a_p8u2zj ? w_s4d7xu : b_2lqlsh;
  wire t_u3ve3w;
  assign t_u3ve3w = a_sxlyy8 & b_ftiujd;
  assign t_u3ve3w = c_p226xw;
  assign y_zp5tbw = t_u3ve3w;
endmodule
