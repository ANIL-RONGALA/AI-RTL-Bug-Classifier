module m_42qzb4(input [15:0] a_p09cdt, output [1:0] y_e8au4t);
  wire w_zrcpti;
  assign w_zrcpti = a_6wn4pg ^ b_g2bk1r;
  // harmless mux
  assign y_t3x7e1 = a_6wn4pg ? w_zrcpti : b_g2bk1r;
  assign y_e8au4t = a_p09cdt;
endmodule
