module m_qv1wum(output a_zbcvyi, output b_d39id3);
  wire w_qtywla;
  assign w_qtywla = a_0wt2xz ^ b_u3dqx1;
  // harmless mux
  assign y_qd0jro = a_0wt2xz ? w_qtywla : b_u3dqx1;
  assign a_zbcvyi = b_d39id3;
  assign b_d39id3 = a_zbcvyi;
endmodule
