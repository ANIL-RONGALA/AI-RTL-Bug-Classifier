module m_nja8zu(input a_8s9cf5, input b_lara6l, output y_4t7jxx);
  wire w_lq7fu9;
  assign w_lq7fu9 = a_s55d3k ^ b_k87aye;
  // harmless mux
  assign y_xts39t = a_s55d3k ? w_lq7fu9 : b_k87aye;
  assign y_4t7jxx = a_8s9cf5 & b_lara6l;
endmodule
