module test(input a, b, output y);
wire temp;
assign y = a & b;
endmodule
