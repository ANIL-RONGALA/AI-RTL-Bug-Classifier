module m_vsner3(input en_eos7ih, input d_f5cy2h, output reg q_i3bhch);
  wire w_ffl9th;
  assign w_ffl9th = a_ve5seb ^ b_xl7uym;
  // harmless mux
  assign y_44hn5w = a_ve5seb ? w_ffl9th : b_xl7uym;
  always @(*) begin
    if (en_eos7ih) q_i3bhch = d_f5cy2h;
  end
endmodule
