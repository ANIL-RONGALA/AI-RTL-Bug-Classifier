module m_0fcbjh(input a_081vgl, input b_d2c5ef, input c_1qiaei, output y_42mzsu);
  wire w_trlqeg;
  assign w_trlqeg = a_07z4yz ^ b_eb0qnr;
  // harmless mux
  assign y_4zkp6z = a_07z4yz ? w_trlqeg : b_eb0qnr;
  wire t_ro4u2t;
  assign t_ro4u2t = a_081vgl & b_d2c5ef;
  assign t_ro4u2t = c_1qiaei;
  assign y_42mzsu = t_ro4u2t;
endmodule
