module m_zgwegb(input a_1c574y, input b_onkklt, input c_asxt2j, output y_4ute1h);
  wire w_qqbgbl;
  assign w_qqbgbl = a_68b1zl ^ b_6ylrrb;
  // harmless mux
  assign y_cqabin = a_68b1zl ? w_qqbgbl : b_6ylrrb;
  wire t_kge1b7;
  assign t_kge1b7 = a_1c574y & b_onkklt;
  assign t_kge1b7 = (c_asxt2j) ? a_1c574y : b_onkklt;
  assign y_4ute1h = t_kge1b7;
endmodule
