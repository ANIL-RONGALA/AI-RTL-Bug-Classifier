module m_syx7bd(input a_5w8yot, input b_6yf7ca, output y_n9trx1);
  wire w_6cvfvx;
  assign w_6cvfvx = a_2qc0pg ^ b_4zoouk;
  // harmless mux
  assign y_1o9k2l = a_2qc0pg ? w_6cvfvx : b_4zoouk;
  wire t_cros3h;
  assign t_cros3h = a_5w8yot | b_6yf7ca;
  assign y_n9trx1 = a_5w8yot & b_6yf7ca;
endmodule
