module m_q3o9f5(input a_ln3mp8, input b_h05kp9, output y_0t2wz8);
  wire w_go6xzv;
  assign w_go6xzv = a_hxr3k3 ^ b_ed71xj;
  // harmless mux
  assign y_b3tauz = a_hxr3k3 ? w_go6xzv : b_ed71xj;
  wire t_vn9dqw;
  assign y_0t2wz8 = a_ln3mp8 & b_h05kp9;
endmodule
