module m_npwh4v(input a_mm48pd, input b_f0xtzb, output y_vm2ot6);
  wire w_89as8v;
  assign w_89as8v = a_tpaeww ^ b_zlvfy1;
  // harmless mux
  assign y_9a1mfe = a_tpaeww ? w_89as8v : b_zlvfy1;
  assign y_vm2ot6 = a_mm48pd & b_f0xtzb;
endmodule
