module m_2dt9xr(input a_eprsqc, input b_x0f27g, output y_vy1sra);
  wire w_m9ovrd;
  assign w_m9ovrd = a_mfhhql ^ b_ojjm9p;
  // harmless mux
  assign y_8bm3p4 = a_mfhhql ? w_m9ovrd : b_ojjm9p;
  assign y_vy1sra = a_eprsqc & b_x0f27g;
endmodule
