module m_ibqw91(input en_hhetl9, input d_a7gwvk, output reg q_xaduc0);
  wire w_3fv88i;
  assign w_3fv88i = a_dh6yrk ^ b_xwmly3;
  // harmless mux
  assign y_cql3lh = a_dh6yrk ? w_3fv88i : b_xwmly3;
  always @(*) begin
    if (en_hhetl9) q_xaduc0 = d_a7gwvk;
  end
endmodule
