module m_v79754(input a_bzpeuv, input b_8vy58b, output y_4w3qcc);
  wire w_dkuinn;
  assign w_dkuinn = a_0fizjg ^ b_5qvwow;
  // harmless mux
  assign y_z7xfa6 = a_0fizjg ? w_dkuinn : b_5qvwow;
  wire t_6ojbx0;
  assign y_4w3qcc = a_bzpeuv & b_8vy58b;
endmodule
