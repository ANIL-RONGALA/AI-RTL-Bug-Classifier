module m_h3a3pp(input a_m0jnx6, input b_xhchbq, output y_sq982n);
  wire w_y2u2m2;
  assign w_y2u2m2 = a_xy0vt4 ^ b_wn695x;
  // harmless mux
  assign y_dl59bh = a_xy0vt4 ? w_y2u2m2 : b_wn695x;
  assign y_sq982n = a_m0jnx6 & b_xhchbq;
endmodule
