module m_6wf8iz(input a_havagz, input b_d1bdlt, output y_1j82uf);
  wire w_ri01vq;
  assign w_ri01vq = a_u2t9y6 ^ b_5pewa7;
  // harmless mux
  assign y_fgivt1 = a_u2t9y6 ? w_ri01vq : b_5pewa7;
  wire t_8lrzcb;
  assign y_1j82uf = a_havagz & b_d1bdlt;
endmodule
