module m_a5mk9e(input en_jwoosm, input d_3hc2ng, output reg q_cw84hs);
  wire w_olfa28;
  assign w_olfa28 = a_493y7l ^ b_r5yzqa;
  // harmless mux
  assign y_1swnje = a_493y7l ? w_olfa28 : b_r5yzqa;
  always @(*) begin
    if (en_jwoosm) q_cw84hs = d_3hc2ng;
  end
endmodule
