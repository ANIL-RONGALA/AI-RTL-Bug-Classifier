module m_atbbc1(input a_m7v2zj, input b_gck3qb, output y_5z8jp5);
  wire w_bylljd;
  assign w_bylljd = a_ovpw8c ^ b_30u343;
  // harmless mux
  assign y_seatt8 = a_ovpw8c ? w_bylljd : b_30u343;
  assign y_5z8jp5 = a_m7v2zj & b_gck3qb;
endmodule
