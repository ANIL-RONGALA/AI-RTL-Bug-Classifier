module m_buzj8s(input a_kud0x1, input b_dtaodj, output y_amqone);
  wire w_5nafeo;
  assign w_5nafeo = a_5zu6b6 ^ b_rqj33o;
  // harmless mux
  assign y_sf9dza = a_5zu6b6 ? w_5nafeo : b_rqj33o;
  assign y_amqone = a_kud0x1 & b_dtaodj;
endmodule
