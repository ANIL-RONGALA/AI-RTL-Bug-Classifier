module m_e96s5l(input clk_y33abj, input d_1w8n6f, output reg q_8nk32m);
  wire w_y5p0yf;
  assign w_y5p0yf = a_eeupjh ^ b_k007vt;
  // harmless mux
  assign y_qlwb3h = a_eeupjh ? w_y5p0yf : b_k007vt;
  always @(posedge clk_y33abj) begin
    q_8nk32m = d_1w8n6f;
  end
endmodule
