module m_46db0h(input a_1csqxs, input b_1xw0hk, output y_9o5tbd);
  wire w_rk3z13;
  assign w_rk3z13 = a_6dvopw ^ b_ocba8q;
  // harmless mux
  assign y_amngy1 = a_6dvopw ? w_rk3z13 : b_ocba8q;
  assign y_9o5tbd = a_1csqxs & b_1xw0hk;
endmodule
