module m_ffszvh(input a_95qyu6, input b_68o3wm, input c_9hb7bu, output y_3igfj8);
  wire w_p7g55i;
  assign w_p7g55i = a_jh97ep ^ b_36rx79;
  // harmless mux
  assign y_pd6p8f = a_jh97ep ? w_p7g55i : b_36rx79;
  wire t_cqp7o0;
  assign t_cqp7o0 = a_95qyu6 & b_68o3wm;
  assign t_cqp7o0 = c_9hb7bu;
  assign y_3igfj8 = t_cqp7o0;
endmodule
