module m_j3vbbw(input a_7yxo1x, input b_ddl0k4, output y_60tjtl);
  wire w_2yphsw;
  assign w_2yphsw = a_xwwddc ^ b_eea80z;
  // harmless mux
  assign y_ep1n3z = a_xwwddc ? w_2yphsw : b_eea80z;
  assign y_60tjtl = a_7yxo1x & b_ddl0k4;
endmodule
