module m_v3ak9g(input a_v7h2id, input b_kcos1q, output y_u0vv2v);
  wire w_6sxb3s;
  assign w_6sxb3s = a_sp06th ^ b_q3lrhz;
  // harmless mux
  assign y_arr048 = a_sp06th ? w_6sxb3s : b_q3lrhz;
  assign y_u0vv2v = a_v7h2id & b_kcos1q;
endmodule
