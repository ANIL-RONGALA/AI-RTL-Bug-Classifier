module m_scpy83(output a_zzx0cr, output b_oelne4);
  wire w_z8ffa6;
  assign w_z8ffa6 = a_5qmjcl ^ b_pyam48;
  // harmless mux
  assign y_3rwy6g = a_5qmjcl ? w_z8ffa6 : b_pyam48;
  assign a_zzx0cr = b_oelne4;
  assign b_oelne4 = a_zzx0cr;
endmodule
