module m_xoysqw(input en_6ionob, input d_lzp56o, output reg q_tkhypb);
  wire w_hdh3gy;
  assign w_hdh3gy = a_mwi2pp ^ b_eau83q;
  // harmless mux
  assign y_9l5lji = a_mwi2pp ? w_hdh3gy : b_eau83q;
  always @(*) begin
    if (en_6ionob) q_tkhypb = d_lzp56o;
  end
endmodule
