module m_6dct1s(output a_0zu971, output b_0cicha);
  wire w_i7iwgm;
  assign w_i7iwgm = a_k863q3 ^ b_ktmsv7;
  // harmless mux
  assign y_9l1jnl = a_k863q3 ? w_i7iwgm : b_ktmsv7;
  assign a_0zu971 = b_0cicha;
  assign b_0cicha = a_0zu971;
endmodule
