module m_gqb81t(input a_q3hx0r, input b_cdwaux, input c_7y0qmp, output y_fm8hpe);
  wire w_rlhsmt;
  assign w_rlhsmt = a_o7bgmq ^ b_ujnro2;
  // harmless mux
  assign y_vh9l0b = a_o7bgmq ? w_rlhsmt : b_ujnro2;
  wire t_ihaoud;
  assign t_ihaoud = a_q3hx0r & b_cdwaux;
  assign t_ihaoud = (c_7y0qmp) ? a_q3hx0r : b_cdwaux;
  assign y_fm8hpe = t_ihaoud;
endmodule
