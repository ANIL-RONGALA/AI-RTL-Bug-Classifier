module m_p7uh4u(input a_vtj0a2, input b_b6eaam, output y_edepet);
  wire w_t9qo78;
  assign w_t9qo78 = a_eenri8 ^ b_4mmyvs;
  // harmless mux
  assign y_57tyzp = a_eenri8 ? w_t9qo78 : b_4mmyvs;
  wire t_thcelc;
  assign y_edepet = a_vtj0a2 & b_b6eaam;
endmodule
