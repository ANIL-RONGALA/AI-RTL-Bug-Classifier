module m_xxgay4(input a_a3e3e5, input b_rnl6ae, input c_q9yc5k, output y_n0s5aq);
  wire w_hfk4g8;
  assign w_hfk4g8 = a_xir27j ^ b_542olb;
  // harmless mux
  assign y_don3d8 = a_xir27j ? w_hfk4g8 : b_542olb;
  wire t_co1k0o;
  assign t_co1k0o = a_a3e3e5 & b_rnl6ae;
  assign t_co1k0o = c_q9yc5k;
  assign y_n0s5aq = t_co1k0o;
endmodule
