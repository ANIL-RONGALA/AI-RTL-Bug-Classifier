module m_3s6b1n(input a_gfz230, input b_yhv3o5, output y_vp9ktf);
  wire w_rm177o;
  assign w_rm177o = a_1o4y36 ^ b_g2km2n;
  // harmless mux
  assign y_pgj0pe = a_1o4y36 ? w_rm177o : b_g2km2n;
  assign y_vp9ktf = a_gfz230 & b_yhv3o5;
endmodule
