module m_vepsne(output a_nkmzgk, output b_sn6im2);
  wire w_1osvqu;
  assign w_1osvqu = a_1du51m ^ b_3006lo;
  // harmless mux
  assign y_w76s7w = a_1du51m ? w_1osvqu : b_3006lo;
  assign a_nkmzgk = b_sn6im2;
  assign b_sn6im2 = a_nkmzgk;
endmodule
