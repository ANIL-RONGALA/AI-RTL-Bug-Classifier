module m_ld6xjn(output a_zmvrmo, output b_w1yney);
  wire w_5ovl8m;
  assign w_5ovl8m = a_r2sxsz ^ b_qk805y;
  // harmless mux
  assign y_92ymhj = a_r2sxsz ? w_5ovl8m : b_qk805y;
  assign a_zmvrmo = b_w1yney;
  assign b_w1yney = a_zmvrmo;
endmodule
