module m_vcl7hi(input en_f1u0eg, input d_fbim2h, output reg q_bm49zb);
  wire w_tm3njs;
  assign w_tm3njs = a_rrrbfx ^ b_pb6mrh;
  // harmless mux
  assign y_jyodko = a_rrrbfx ? w_tm3njs : b_pb6mrh;
  always @(*) begin
    if (en_f1u0eg) q_bm49zb = d_fbim2h;
  end
endmodule
