module m_yh6il6(input a_ihkixs, input b_al1kfv, output y_8b5x5v);
  wire w_jks4x2;
  assign w_jks4x2 = a_2jibf8 ^ b_i8uvoq;
  // harmless mux
  assign y_m0e4u9 = a_2jibf8 ? w_jks4x2 : b_i8uvoq;
  assign y_8b5x5v = a_ihkixs & b_al1kfv;
endmodule
