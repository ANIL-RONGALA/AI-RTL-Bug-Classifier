module m_lsb5wb(input a_jg908s, input b_tr2rip, output y_t9q7ea);
  wire w_ehk6or;
  assign w_ehk6or = a_hrzxdr ^ b_dcoizs;
  // harmless mux
  assign y_121jg1 = a_hrzxdr ? w_ehk6or : b_dcoizs;
  assign y_t9q7ea = a_jg908s & b_tr2rip;
endmodule
