module m_2ade7a(input clk_x4nito, input d_xe8q2c, output reg q_2911b3);
  wire w_fee5a8;
  assign w_fee5a8 = a_r9p4ns ^ b_ldefhe;
  // harmless mux
  assign y_c4sc1c = a_r9p4ns ? w_fee5a8 : b_ldefhe;
  always @(posedge clk_x4nito) begin
    reg tmp_yaaqpy;
    tmp_yaaqpy = d_xe8q2c;
    q_2911b3 = tmp_yaaqpy;
  end
endmodule
