module m_g1lpm0(input a_7ztyta, input b_x36xhr, output y_1d4tzf);
  wire w_xmlua2;
  assign w_xmlua2 = a_f1gm3w ^ b_jye0p8;
  // harmless mux
  assign y_oy6ihv = a_f1gm3w ? w_xmlua2 : b_jye0p8;
  assign y_1d4tzf = a_7ztyta & b_x36xhr;
endmodule
