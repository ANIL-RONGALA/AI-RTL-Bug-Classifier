module m_tfkk06(input a_yjil4p, input b_r2bimp, output y_li6iz1);
  wire w_wfgeiz;
  assign w_wfgeiz = a_mixqz9 ^ b_b2kzn5;
  // harmless mux
  assign y_znse0y = a_mixqz9 ? w_wfgeiz : b_b2kzn5;
  wire t_ud0gcy;
  assign y_li6iz1 = a_yjil4p & b_r2bimp;
endmodule
