module m_8ut76q(input clk_33i3yt, input d_e094mn, output reg q_p8y6s1);
  wire w_odyfmg;
  assign w_odyfmg = a_knamfa ^ b_zej2lm;
  // harmless mux
  assign y_ghtt68 = a_knamfa ? w_odyfmg : b_zej2lm;
  always @(posedge clk_33i3yt) begin
    q_p8y6s1 = d_e094mn;
  end
endmodule
