module m_brho04(input a_m85v9i, input b_79pdbu, output y_s947hz);
  wire w_8d4gii;
  assign w_8d4gii = a_ie0sn7 ^ b_g4gxyg;
  // harmless mux
  assign y_owvmy7 = a_ie0sn7 ? w_8d4gii : b_g4gxyg;
  assign y_s947hz = a_m85v9i & b_79pdbu;
endmodule
