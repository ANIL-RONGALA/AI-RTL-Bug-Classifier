module m_3l39g0(input clk_qemxxl, input d_cxjw5l, output reg q_arzpih);
  wire w_dx9ror;
  assign w_dx9ror = a_1fy1uf ^ b_vh27aj;
  // harmless mux
  assign y_mods04 = a_1fy1uf ? w_dx9ror : b_vh27aj;
  always @(posedge clk_qemxxl) begin
    reg tmp_eivz1a;
    tmp_eivz1a = d_cxjw5l;
    q_arzpih = tmp_eivz1a;
  end
endmodule
