module m_5m1sel(input a_hnjmg0, input b_u1wqhh, output y_7s88nc);
  wire w_llfvp7;
  assign w_llfvp7 = a_67bvad ^ b_xqhuoa;
  // harmless mux
  assign y_vaolb4 = a_67bvad ? w_llfvp7 : b_xqhuoa;
  assign y_7s88nc = a_hnjmg0 & b_u1wqhh;
endmodule
