module m_86yzv7(input a_qy9pl2, input b_31z8wm, output y_ajwu9a);
  wire w_u75qfh;
  assign w_u75qfh = a_x6uiti ^ b_wvpqjn;
  // harmless mux
  assign y_p73afh = a_x6uiti ? w_u75qfh : b_wvpqjn;
  assign y_ajwu9a = a_qy9pl2 & b_31z8wm;
endmodule
