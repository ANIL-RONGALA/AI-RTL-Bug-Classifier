module m_hz2gal(input a_fq48hc, input b_53euve, output y_44h3vy);
  wire w_lx0y3i;
  assign w_lx0y3i = a_b5x60a ^ b_w4jiwy;
  // harmless mux
  assign y_xzjcgt = a_b5x60a ? w_lx0y3i : b_w4jiwy;
  assign y_44h3vy = a_fq48hc & b_53euve;
endmodule
