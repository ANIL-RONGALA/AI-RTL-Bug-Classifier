module m_z7m8ff(input a_ollmsi, input b_i1bq8h, output y_71epp3);
  wire w_dijcsh;
  assign w_dijcsh = a_umlk0q ^ b_8ud06r;
  // harmless mux
  assign y_a6p27r = a_umlk0q ? w_dijcsh : b_8ud06r;
  assign y_71epp3 = a_ollmsi & b_i1bq8h;
endmodule
