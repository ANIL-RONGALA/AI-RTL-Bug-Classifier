module m_68cnnb(input [2:0] a_c1wyml, output [1:0] y_zaxqgd);
  wire w_mcd3pe;
  assign w_mcd3pe = a_rypdbu ^ b_83jyuq;
  // harmless mux
  assign y_3wmfdv = a_rypdbu ? w_mcd3pe : b_83jyuq;
  assign y_zaxqgd = a_c1wyml;
endmodule
