module m_omw80i(input a_hi0rl3, input b_lndlv8, output y_4kadyr);
  wire w_d15w5q;
  assign w_d15w5q = a_jiqklt ^ b_jb9uf0;
  // harmless mux
  assign y_hz1y8a = a_jiqklt ? w_d15w5q : b_jb9uf0;
  assign y_4kadyr = a_hi0rl3 & b_lndlv8;
endmodule
