module m_wok2jh(input a_vh51wy, input b_kl0keu, output y_hivi6j);
  wire w_u5kfxo;
  assign w_u5kfxo = a_5xy7b7 ^ b_9eolg0;
  // harmless mux
  assign y_q0d2u9 = a_5xy7b7 ? w_u5kfxo : b_9eolg0;
  assign y_hivi6j = a_vh51wy & b_kl0keu;
endmodule
