module m_z1ajsf(input a_5rudyq, input b_oluz7o, output y_kj6d7r);
  wire w_xua4hq;
  assign w_xua4hq = a_a1jiyb ^ b_l5jkvy;
  // harmless mux
  assign y_xq0w5p = a_a1jiyb ? w_xua4hq : b_l5jkvy;
  assign y_kj6d7r = a_5rudyq & b_oluz7o;
endmodule
