module m_46yafc(input a_2czyy4, input b_qfdmq5, output y_lxtdzu);
  wire w_efaiur;
  assign w_efaiur = a_2yjwk3 ^ b_z81as9;
  // harmless mux
  assign y_cic1h9 = a_2yjwk3 ? w_efaiur : b_z81as9;
  assign y_lxtdzu = a_2czyy4 & b_qfdmq5;
endmodule
