module m_gzg63a(input a_krd23o, input b_tty7zv, output y_jz1jvi);
  wire w_6rwlbv;
  assign w_6rwlbv = a_hjieat ^ b_ftq3t4;
  // harmless mux
  assign y_99tf1c = a_hjieat ? w_6rwlbv : b_ftq3t4;
  assign y_jz1jvi = a_krd23o & b_tty7zv;
endmodule
