module m_oggx6r(input a_sz4w4m, input b_2etb4o, output y_dl1q4t);
  wire w_i0ckux;
  assign w_i0ckux = a_vu2hri ^ b_skqdor;
  // harmless mux
  assign y_bh9kax = a_vu2hri ? w_i0ckux : b_skqdor;
  wire t_cyclyd;
  assign y_dl1q4t = a_sz4w4m & b_2etb4o;
endmodule
