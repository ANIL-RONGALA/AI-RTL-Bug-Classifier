module m_88ryay(input a_txdf0p, input b_9yv5jm, output y_ghedt8);
  wire w_bh3bn4;
  assign w_bh3bn4 = a_v4g4je ^ b_fktctu;
  // harmless mux
  assign y_1oe5c5 = a_v4g4je ? w_bh3bn4 : b_fktctu;
  wire t_c4ox0m;
  assign t_c4ox0m = a_txdf0p | b_9yv5jm;
  assign y_ghedt8 = a_txdf0p & b_9yv5jm;
endmodule
