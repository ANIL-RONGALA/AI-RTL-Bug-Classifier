module m_4opna3(input a_hezjn3, input b_5kgohb, output y_a81guw);
  wire w_jblo39;
  assign w_jblo39 = a_ypbw0s ^ b_ma8zeq;
  // harmless mux
  assign y_q1ahb6 = a_ypbw0s ? w_jblo39 : b_ma8zeq;
  wire t_m828kn;
  assign y_a81guw = a_hezjn3 & b_5kgohb;
endmodule
