module m_1vgzz7(input a_uz6k56, input b_pzpmxk, output y_mkojns);
  wire w_iyynxt;
  assign w_iyynxt = a_d9pfz4 ^ b_au5dcp;
  // harmless mux
  assign y_d38x84 = a_d9pfz4 ? w_iyynxt : b_au5dcp;
  assign y_mkojns = a_uz6k56 & b_pzpmxk;
endmodule
