module m_cu2m83(input a_10hcjm, input b_s3fs3r, output y_0cmlt1);
  wire w_mb5jl4;
  assign w_mb5jl4 = a_rkdv9c ^ b_uq3cf3;
  // harmless mux
  assign y_v971bj = a_rkdv9c ? w_mb5jl4 : b_uq3cf3;
  wire t_mn1pfk;
  assign t_mn1pfk = a_10hcjm | b_s3fs3r;
  assign y_0cmlt1 = a_10hcjm & b_s3fs3r;
endmodule
