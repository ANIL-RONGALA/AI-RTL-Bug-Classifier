module m_fs1lea(input a_16yqp7, input b_llpri3, output y_4s85fb);
  wire w_f2zcce;
  assign w_f2zcce = a_w1rj3i ^ b_zhr6ue;
  // harmless mux
  assign y_jpqxmp = a_w1rj3i ? w_f2zcce : b_zhr6ue;
  assign y_4s85fb = a_16yqp7 & b_llpri3;
endmodule
