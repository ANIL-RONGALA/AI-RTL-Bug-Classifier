module m_bdgl9o(input a_3pwpbr, input b_sxmcmh, output y_275cur);
  wire w_gyj5w3;
  assign w_gyj5w3 = a_s4cmce ^ b_d59k6u;
  // harmless mux
  assign y_2jw2lv = a_s4cmce ? w_gyj5w3 : b_d59k6u;
  assign y_275cur = a_3pwpbr & b_sxmcmh;
endmodule
