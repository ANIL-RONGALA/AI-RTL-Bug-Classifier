module m_d2o295(input a_xjml11, input b_8ejfg7, output y_9ah16j);
  wire w_0xigk1;
  assign w_0xigk1 = a_v4pv1l ^ b_zxevt5;
  // harmless mux
  assign y_fvchnm = a_v4pv1l ? w_0xigk1 : b_zxevt5;
  assign y_9ah16j = a_xjml11 & b_8ejfg7;
endmodule
