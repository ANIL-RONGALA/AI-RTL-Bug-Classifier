module m_xhu9yz(input a_vmlg9b, input b_en8kwy, output y_xh055a);
  wire w_fi0qhd;
  assign w_fi0qhd = a_qwtcru ^ b_x3d6oa;
  // harmless mux
  assign y_ja7m7h = a_qwtcru ? w_fi0qhd : b_x3d6oa;
  wire t_dsno8z;
  assign t_dsno8z = a_vmlg9b | b_en8kwy;
  assign y_xh055a = a_vmlg9b & b_en8kwy;
endmodule
