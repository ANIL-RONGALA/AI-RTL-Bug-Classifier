module m_yfeevn(input a_z8xu18, input b_ubjv6j, output y_gfcc9o);
  wire w_q4qf97;
  assign w_q4qf97 = a_42m8v1 ^ b_of8ex6;
  // harmless mux
  assign y_59m87a = a_42m8v1 ? w_q4qf97 : b_of8ex6;
  assign y_gfcc9o = a_z8xu18 & b_ubjv6j;
endmodule
