module m_2purru(input [3:0] a_r37q32, output [2:0] y_6t956b);
  wire w_5on2dh;
  assign w_5on2dh = a_1mybg1 ^ b_zq27ve;
  // harmless mux
  assign y_em5pwu = a_1mybg1 ? w_5on2dh : b_zq27ve;
  assign y_6t956b = a_r37q32;
endmodule
