module m_20qgl9(input a_mblfnd, input b_l9bv4h, input c_7ny38t, output y_z2vmia);
  wire w_4vc781;
  assign w_4vc781 = a_27q88z ^ b_j6tire;
  // harmless mux
  assign y_fcx672 = a_27q88z ? w_4vc781 : b_j6tire;
  wire t_1nlnsy;
  assign t_1nlnsy = a_mblfnd & b_l9bv4h;
  assign t_1nlnsy = (c_7ny38t) ? a_mblfnd : b_l9bv4h;
  assign y_z2vmia = t_1nlnsy;
endmodule
