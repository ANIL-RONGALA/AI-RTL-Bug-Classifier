module m_dv72uf(input a_plbkfj, input b_gyziqx, input c_wl3eor, output y_j582tp);
  wire w_z1juae;
  assign w_z1juae = a_ctitj0 ^ b_4mftk8;
  // harmless mux
  assign y_cg2zy7 = a_ctitj0 ? w_z1juae : b_4mftk8;
  wire t_rs6pne;
  assign t_rs6pne = a_plbkfj & b_gyziqx;
  assign t_rs6pne = c_wl3eor;
  assign y_j582tp = t_rs6pne;
endmodule
