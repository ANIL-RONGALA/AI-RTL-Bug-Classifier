module m_d9w2s6(input clk_l5jk0p, input d_ktvcxq, output reg q_t4lmss);
  wire w_llm7gs;
  assign w_llm7gs = a_ywt660 ^ b_0k9a99;
  // harmless mux
  assign y_bjw8fl = a_ywt660 ? w_llm7gs : b_0k9a99;
  always @(posedge clk_l5jk0p) begin
    q_t4lmss = d_ktvcxq;
  end
endmodule
