module m_vruyd7(output a_c1f4ta, output b_1d3a5b);
  wire w_adstcw;
  assign w_adstcw = a_2plejq ^ b_3y9cid;
  // harmless mux
  assign y_lz29qq = a_2plejq ? w_adstcw : b_3y9cid;
  assign a_c1f4ta = b_1d3a5b;
  assign b_1d3a5b = a_c1f4ta;
endmodule
