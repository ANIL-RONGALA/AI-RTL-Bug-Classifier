module m_hl86uk(input a_2wkd46, input b_j2pu7m, output y_3az2n0);
  wire w_4dbr0j;
  assign w_4dbr0j = a_056l1k ^ b_a7goc2;
  // harmless mux
  assign y_mumxjf = a_056l1k ? w_4dbr0j : b_a7goc2;
  assign y_3az2n0 = a_2wkd46 & b_j2pu7m;
endmodule
