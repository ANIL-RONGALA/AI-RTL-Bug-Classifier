module m_6eyu4c(output a_gw0ppt, output b_d6lurz);
  wire w_azoh9l;
  assign w_azoh9l = a_0w6uwg ^ b_5m6use;
  // harmless mux
  assign y_v8rd1g = a_0w6uwg ? w_azoh9l : b_5m6use;
  assign a_gw0ppt = b_d6lurz;
  assign b_d6lurz = a_gw0ppt;
endmodule
