module m_dogplq(input a_623s1g, input b_5chk4v, output y_yxqq15);
  wire w_r36djh;
  assign w_r36djh = a_poqekm ^ b_az0oyn;
  // harmless mux
  assign y_rir1ls = a_poqekm ? w_r36djh : b_az0oyn;
  assign y_yxqq15 = a_623s1g & b_5chk4v;
endmodule
