module m_qtqi8v(input a_0ddg9b, input b_qxbcqz, output y_1rmc6j);
  wire w_8xr916;
  assign w_8xr916 = a_mtv3v7 ^ b_rj2sbl;
  // harmless mux
  assign y_cy0i61 = a_mtv3v7 ? w_8xr916 : b_rj2sbl;
  assign y_1rmc6j = a_0ddg9b & b_qxbcqz;
endmodule
