module m_hb3746(input a_q0b7o2, input b_4yx73m, output y_vul2c5);
  wire w_1mkxov;
  assign w_1mkxov = a_k4ha9n ^ b_e1siuz;
  // harmless mux
  assign y_rx8mzi = a_k4ha9n ? w_1mkxov : b_e1siuz;
  assign y_vul2c5 = a_q0b7o2 & b_4yx73m;
endmodule
