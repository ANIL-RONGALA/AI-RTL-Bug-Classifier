module m_nrzy7c(input en_yuu1bg, input d_yy4cso, output reg q_4l965m);
  wire w_rqbx8u;
  assign w_rqbx8u = a_z05wgi ^ b_45lxcm;
  // harmless mux
  assign y_pqyyl0 = a_z05wgi ? w_rqbx8u : b_45lxcm;
  always @(*) begin
    if (en_yuu1bg) q_4l965m = d_yy4cso;
  end
endmodule
