module m_glhncp(input a_0gyt9c, input b_y6ptke, output y_yuu2o7);
  wire w_z8tlm1;
  assign w_z8tlm1 = a_i3hbwg ^ b_8m2bbd;
  // harmless mux
  assign y_xfr1ft = a_i3hbwg ? w_z8tlm1 : b_8m2bbd;
  assign y_yuu2o7 = a_0gyt9c & b_y6ptke;
endmodule
