module m_8s4b3c(input en_zg5a6p, input d_32mcuo, output reg q_5v9pvl);
  wire w_gfgqwf;
  assign w_gfgqwf = a_myviio ^ b_p4year;
  // harmless mux
  assign y_97segd = a_myviio ? w_gfgqwf : b_p4year;
  always @(*) begin
    if (en_zg5a6p) q_5v9pvl = d_32mcuo;
  end
endmodule
